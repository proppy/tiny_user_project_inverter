* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output12_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput10 net10 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput9 net9 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput11 net11 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput12 net12 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output10_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net13 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_007_ net6 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__004__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput14 net14 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_006_ net7 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__007__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput15 net15 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_005_ net8 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput16 net16 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_004_ net1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_003_ net2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_002_ net3 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_001_ net4 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_180 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_000_ net5 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_170 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_181 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_160 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_182 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_171 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_150 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_161 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_183 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_172 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_151 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_133_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_140 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_162 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_184 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_173 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_90 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_130 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_141 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_174 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_163 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_152 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_91 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput5 io_in[14] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_80 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__002__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_131 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_120 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_142 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_175 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_164 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_153 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__005__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput6 io_in[15] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_81 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_70 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_92 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_121 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_110 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_132 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_143 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_165 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_154 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_176 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_93 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_71 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput7 io_in[8] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_82 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_60 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_122 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_111 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_100 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_133 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_166 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_144 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_155 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_177 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_50 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_72 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 io_in[9] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_61 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_83 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_94 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_101 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_112 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_123 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_134 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_145 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_156 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_167 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_178 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_40 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_84 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_62 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_51 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_73 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_95 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_180_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_124 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_102 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_113 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_146 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_135 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_157 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_168 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_179 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_41 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_30 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_74 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_63 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_96 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_85 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_103 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_114 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_147 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_125 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_136 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_169 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_158 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_31 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_20 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_64 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_53 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_75 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_42 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_86 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_97 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_104 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_115 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_126 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_137 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_148 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_159 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_21 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_32 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_43 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_54 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_65 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_76 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_98 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_87 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_185_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_92_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_92_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_105 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_116 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_127 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_138 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_149 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_22 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_44 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_33 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_55 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_66 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_77 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_88 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_99 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_180_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_106 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_139 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_117 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_128 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_23 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_34 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_45 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_56 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_67 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_78 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_89 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_118 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_129 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_107 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_24 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_35 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_57 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_46 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_68 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_79 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_195_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_119 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_108 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_47 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_25 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_36 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_69 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_58 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_195_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_109 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__000__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_26 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_37 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_48 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_59 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__003__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_38 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_27 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_49 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__006__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_17 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_39 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_28 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_29 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_18 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_19 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

